module backend

pub const (
	i_am_being_used = 420
)

pub fn init() {
	println("[BACKEND] TODO")
}