module enums

pub const (
	clip_part = 1
	clip_all  = 2
)

pub const (
	command_jump = 1
	command_clip = 2
	command_rect = 3
	command_text = 4
	command_icon = 5
	command_max  = 6
)

pub const (
	color_text        = 0
	color_border      = 1
	color_windowbg    = 2
	color_titlebg     = 3
	color_titletext   = 4
	color_panelbg     = 5
	color_button      = 6
	color_buttonhover = 7
	color_buttonfocus = 8
	color_base        = 9
	color_basehover   = 10
	color_basefocus   = 11
	color_scrollbase  = 12
	color_scrollthumb = 13
	color_max         = 14
)
