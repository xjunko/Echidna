module common

pub enum MouseButton {
	left
	middle
	right
}
