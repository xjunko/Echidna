module vector

// Shortcuts, i dont really use this doe
pub type Vector2f = Vector2<f64>
pub type Vector2i = Vector2<int>